`include "config.svh"

module lab_top
# (
    parameter  clk_mhz       = 50,
               w_key         = 4,
               w_sw          = 8,
               w_led         = 8,
               w_digit       = 8,
               w_gpio        = 100,

               screen_width  = 640,
               screen_height = 480,

               w_red         = 4,
               w_green       = 4,
               w_blue        = 4,

               w_x           = $clog2 ( screen_width  ),
               w_y           = $clog2 ( screen_height )
)
(
    input                        clk,
    input                        slow_clk,
    input                        rst,

    // Keys, switches, LEDs

    input        [w_key   - 1:0] key,
    input        [w_sw    - 1:0] sw,
    output logic [w_led   - 1:0] led,

    // A dynamic seven-segment display

    output logic [          7:0] abcdefgh,
    output logic [w_digit - 1:0] digit,

    // Graphics

    input        [w_x     - 1:0] x,
    input        [w_y     - 1:0] y,

    output logic [w_red   - 1:0] red,
    output logic [w_green - 1:0] green,
    output logic [w_blue  - 1:0] blue,

    // Microphone, sound output and UART

    input        [         23:0] mic,
    output       [         15:0] sound,

    input                        uart_rx,
    output                       uart_tx,

    // General-purpose Input/Output

    inout        [w_gpio  - 1:0] gpio
);

    //------------------------------------------------------------------------

    // assign led        = '0;
    // assign abcdefgh   = '0;
    // assign digit      = '0;
       assign red        = '0;
       assign green      = '0;
       assign blue       = '0;
       assign sound      = '0;
       assign uart_tx    = '1;

    //------------------------------------------------------------------------

    logic [31:0] cnt;

    always_ff @ (posedge clk or posedge rst)
        if (rst)
            cnt <= '0;
        else
            cnt <= cnt + 1'd1;

    // wire enable = (cnt [24:0] == '0);
    wire enable;

    //------------------------------------------------------------------------

    logic [w_digit:0] shift_reg;

    always_ff @ (posedge clk or posedge rst)
      if (rst)
        shift_reg <= w_digit' (1);
      else if (enable)
        shift_reg <= { shift_reg [0], shift_reg [w_digit - 1:1] };

    assign led[8:0] = (w_led)' (shift_reg);

    //------------------------------------------------------------------------

    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d--  h

    typedef enum bit [7:0]
    {
        F     = 8'b1000_1110,
        P     = 8'b1100_1110,
        G     = 8'b1011_1100,
        A     = 8'b1110_1110,
        space = 8'b0000_0000
    }
    seven_seg_encoding_e;

    // seven_seg_encoding_e letter;
    wire [7:0] letter;

    // always_comb
    //   case (4' (shift_reg))
    //   4'b1000: letter = F;
    //   4'b0100: letter = P;
    //   4'b0010: letter = G;
    //   4'b0001: letter = A;
    //   default: letter = space;
    //   endcase

    assign abcdefgh = letter;
    assign digit    = shift_reg;

    // Recieve with laser
    wire uart_in = ~ gpio[30];

    uart_rx #(
        .CLK_FREQ  (  50000000 ), // clk frequency, Unit : Hz
        .BAUD_RATE (  1200     ), // Unit : Hz
        .PARITY    (  "NONE"   ), // "NONE", "ODD", or "EVEN"
        .FIFO_EA   (  3        ) // 0:no fifo   1,2:depth=4   3:depth=8   4:depth=16  ...  10:depth=1024   11:depth=2048  ...
    ) (
        .rstn       ( ~rst ),
        .clk        ( clk  ),

        .i_uart_rx  ( uart_in ),

        .o_tready   ( '1     ),
        .o_tvalid   ( enable ),
        .o_tdata    ( letter ),
        .o_overflow (  )
    );

    assign led[9] = uart_in;

endmodule
